
package tb_pkg;

`include "uvm_macros.svh"

import i2c_vip_pkg::*;
import spi_vip_pkg::*;
import axi4stream_vip_pkg::*;
import axis_master_0_pkg::*;
import axis_slave_0_pkg::*;
import axi4stream_uvm_pkg::*;
import axis_i2c_master_pkg::*;
import uvm_pkg::*;

`include "tests/basic_test.svh"

endpackage