module tb_top_deserialized(

    );

    spi_intf spi_if();
endmodule
