package axi4stream_uvm_pkg;

`include "uvm_macros.svh"
import uvm_pkg::*;
import axi4stream_vip_pkg::*;
import generic_components_pkg::*;

`include "axi4stream_uvm_transaction.svh"
`include "axi4stream_uvm_mst_agent.svh"
`include "axi4stream_uvm_slv_agent.svh"
`include "byteq_to_axi4stream.svh"

endpackage