package spi_vip_pkg;

`include "uvm_macros.svh"
import uvm_pkg::*;

`include "spi_item.svh"
`include "spi_monitor.svh"
`include "spi_mst_driver.svh"

endpackage