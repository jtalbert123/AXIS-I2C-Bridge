

package generic_components_pkg;

`include "uvm_macros.svh"
import uvm_pkg::*;

`include "generic_listener.svh"
`include "byteq.svh"

endpackage